module neurona1()